module static_not_taken (

	output logic br_predict
	
);

assign br_predict = 1'b0;

endmodule : static_not_taken